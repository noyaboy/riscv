
module Icache #(
            parameter ADDR_WIDTH = 8,
            parameter ADDR_NUM = 256
        ) (
            input clk,
            input rst_n,
            input wen,
            input pc_running,
            input [7:0] boot_addr,
            input [31:0] pc, 
            input [32-1:0] wdata,
            output reg [32-1: 0] rdata
        );
/*
reg [32-1: 0] mem [256-1: 0];
reg [32-1: 0] mem_n [256-1: 0];
integer i;

always @ (posedge clk) 
    if (~rst_n) begin
        for(i = 0; i < ADDR_NUM; i = i + 1) mem[i] <= 0;
    end
    else begin
        for(i = 0; i < ADDR_NUM; i = i + 1) mem[i] <= mem_n[i];
    end

always@* 
    rdata = mem[addr];

always @(*) begin
	for(i = 0; i < ADDR_NUM; i = i + 1) begin
		mem_n[i] = (wen && (i == addr)) ? wdata : mem[i];
	end
end
*/
wire [ADDR_WIDTH-1: 0] addr;
assign addr = pc_running ? pc[ADDR_WIDTH + 1: 2] : boot_addr;

reg [32-1: 0] mem0;
    reg [32-1: 0] mem1;
    reg [32-1: 0] mem2;
    reg [32-1: 0] mem3;
    reg [32-1: 0] mem4;
    reg [32-1: 0] mem5;
    reg [32-1: 0] mem6;
    reg [32-1: 0] mem7;
    reg [32-1: 0] mem8;
    reg [32-1: 0] mem9;
    reg [32-1: 0] mem10;
    reg [32-1: 0] mem11;
    reg [32-1: 0] mem12;
    reg [32-1: 0] mem13;
    reg [32-1: 0] mem14;
    reg [32-1: 0] mem15;
    reg [32-1: 0] mem16;
    reg [32-1: 0] mem17;
    reg [32-1: 0] mem18;
    reg [32-1: 0] mem19;
    reg [32-1: 0] mem20;
    reg [32-1: 0] mem21;
    reg [32-1: 0] mem22;
    reg [32-1: 0] mem23;
    reg [32-1: 0] mem24;
    reg [32-1: 0] mem25;
    reg [32-1: 0] mem26;
    reg [32-1: 0] mem27;
    reg [32-1: 0] mem28;
    reg [32-1: 0] mem29;
    reg [32-1: 0] mem30;
    reg [32-1: 0] mem31;
    reg [32-1: 0] mem32;
    reg [32-1: 0] mem33;
    reg [32-1: 0] mem34;
    reg [32-1: 0] mem35;
    reg [32-1: 0] mem36;
    reg [32-1: 0] mem37;
    reg [32-1: 0] mem38;
    reg [32-1: 0] mem39;
    reg [32-1: 0] mem40;
    reg [32-1: 0] mem41;
    reg [32-1: 0] mem42;
    reg [32-1: 0] mem43;
    reg [32-1: 0] mem44;
    reg [32-1: 0] mem45;
    reg [32-1: 0] mem46;
    reg [32-1: 0] mem47;
    reg [32-1: 0] mem48;
    reg [32-1: 0] mem49;
    reg [32-1: 0] mem50;
    reg [32-1: 0] mem51;
    reg [32-1: 0] mem52;
    reg [32-1: 0] mem53;
    reg [32-1: 0] mem54;
    reg [32-1: 0] mem55;
    reg [32-1: 0] mem56;
    reg [32-1: 0] mem57;
    reg [32-1: 0] mem58;
    reg [32-1: 0] mem59;
    reg [32-1: 0] mem60;
    reg [32-1: 0] mem61;
    reg [32-1: 0] mem62;
    reg [32-1: 0] mem63;
    reg [32-1: 0] mem64;
    reg [32-1: 0] mem65;
    reg [32-1: 0] mem66;
    reg [32-1: 0] mem67;
    reg [32-1: 0] mem68;
    reg [32-1: 0] mem69;
    reg [32-1: 0] mem70;
    reg [32-1: 0] mem71;
    reg [32-1: 0] mem72;
    reg [32-1: 0] mem73;
    reg [32-1: 0] mem74;
    reg [32-1: 0] mem75;
    reg [32-1: 0] mem76;
    reg [32-1: 0] mem77;
    reg [32-1: 0] mem78;
    reg [32-1: 0] mem79;
    reg [32-1: 0] mem80;
    reg [32-1: 0] mem81;
    reg [32-1: 0] mem82;
    reg [32-1: 0] mem83;
    reg [32-1: 0] mem84;
    reg [32-1: 0] mem85;
    reg [32-1: 0] mem86;
    reg [32-1: 0] mem87;
    reg [32-1: 0] mem88;
    reg [32-1: 0] mem89;
    reg [32-1: 0] mem90;
    reg [32-1: 0] mem91;
    reg [32-1: 0] mem92;
    reg [32-1: 0] mem93;
    reg [32-1: 0] mem94;
    reg [32-1: 0] mem95;
    reg [32-1: 0] mem96;
    reg [32-1: 0] mem97;
    reg [32-1: 0] mem98;
    reg [32-1: 0] mem99;
    reg [32-1: 0] mem100;
    reg [32-1: 0] mem101;
    reg [32-1: 0] mem102;
    reg [32-1: 0] mem103;
    reg [32-1: 0] mem104;
    reg [32-1: 0] mem105;
    reg [32-1: 0] mem106;
    reg [32-1: 0] mem107;
    reg [32-1: 0] mem108;
    reg [32-1: 0] mem109;
    reg [32-1: 0] mem110;
    reg [32-1: 0] mem111;
    reg [32-1: 0] mem112;
    reg [32-1: 0] mem113;
    reg [32-1: 0] mem114;
    reg [32-1: 0] mem115;
    reg [32-1: 0] mem116;
    reg [32-1: 0] mem117;
    reg [32-1: 0] mem118;
    reg [32-1: 0] mem119;
    reg [32-1: 0] mem120;
    reg [32-1: 0] mem121;
    reg [32-1: 0] mem122;
    reg [32-1: 0] mem123;
    reg [32-1: 0] mem124;
    reg [32-1: 0] mem125;
    reg [32-1: 0] mem126;
    reg [32-1: 0] mem127;
    reg [32-1: 0] mem128;
    reg [32-1: 0] mem129;
    reg [32-1: 0] mem130;
    reg [32-1: 0] mem131;
    reg [32-1: 0] mem132;
    reg [32-1: 0] mem133;
    reg [32-1: 0] mem134;
    reg [32-1: 0] mem135;
    reg [32-1: 0] mem136;
    reg [32-1: 0] mem137;
    reg [32-1: 0] mem138;
    reg [32-1: 0] mem139;
    reg [32-1: 0] mem140;
    reg [32-1: 0] mem141;
    reg [32-1: 0] mem142;
    reg [32-1: 0] mem143;
    reg [32-1: 0] mem144;
    reg [32-1: 0] mem145;
    reg [32-1: 0] mem146;
    reg [32-1: 0] mem147;
    reg [32-1: 0] mem148;
    reg [32-1: 0] mem149;
    reg [32-1: 0] mem150;
    reg [32-1: 0] mem151;
    reg [32-1: 0] mem152;
    reg [32-1: 0] mem153;
    reg [32-1: 0] mem154;
    reg [32-1: 0] mem155;
    reg [32-1: 0] mem156;
    reg [32-1: 0] mem157;
    reg [32-1: 0] mem158;
    reg [32-1: 0] mem159;
    reg [32-1: 0] mem160;
    reg [32-1: 0] mem161;
    reg [32-1: 0] mem162;
    reg [32-1: 0] mem163;
    reg [32-1: 0] mem164;
    reg [32-1: 0] mem165;
    reg [32-1: 0] mem166;
    reg [32-1: 0] mem167;
    reg [32-1: 0] mem168;
    reg [32-1: 0] mem169;
    reg [32-1: 0] mem170;
    reg [32-1: 0] mem171;
    reg [32-1: 0] mem172;
    reg [32-1: 0] mem173;
    reg [32-1: 0] mem174;
    reg [32-1: 0] mem175;
    reg [32-1: 0] mem176;
    reg [32-1: 0] mem177;
    reg [32-1: 0] mem178;
    reg [32-1: 0] mem179;
    reg [32-1: 0] mem180;
    reg [32-1: 0] mem181;
    reg [32-1: 0] mem182;
    reg [32-1: 0] mem183;
    reg [32-1: 0] mem184;
    reg [32-1: 0] mem185;
    reg [32-1: 0] mem186;
    reg [32-1: 0] mem187;
    reg [32-1: 0] mem188;
    reg [32-1: 0] mem189;
    reg [32-1: 0] mem190;
    reg [32-1: 0] mem191;
    reg [32-1: 0] mem192;
    reg [32-1: 0] mem193;
    reg [32-1: 0] mem194;
    reg [32-1: 0] mem195;
    reg [32-1: 0] mem196;
    reg [32-1: 0] mem197;
    reg [32-1: 0] mem198;
    reg [32-1: 0] mem199;
    reg [32-1: 0] mem200;
    reg [32-1: 0] mem201;
    reg [32-1: 0] mem202;
    reg [32-1: 0] mem203;
    reg [32-1: 0] mem204;
    reg [32-1: 0] mem205;
    reg [32-1: 0] mem206;
    reg [32-1: 0] mem207;
    reg [32-1: 0] mem208;
    reg [32-1: 0] mem209;
    reg [32-1: 0] mem210;
    reg [32-1: 0] mem211;
    reg [32-1: 0] mem212;
    reg [32-1: 0] mem213;
    reg [32-1: 0] mem214;
    reg [32-1: 0] mem215;
    reg [32-1: 0] mem216;
    reg [32-1: 0] mem217;
    reg [32-1: 0] mem218;
    reg [32-1: 0] mem219;
    reg [32-1: 0] mem220;
    reg [32-1: 0] mem221;
    reg [32-1: 0] mem222;
    reg [32-1: 0] mem223;
    reg [32-1: 0] mem224;
    reg [32-1: 0] mem225;
    reg [32-1: 0] mem226;
    reg [32-1: 0] mem227;
    reg [32-1: 0] mem228;
    reg [32-1: 0] mem229;
    reg [32-1: 0] mem230;
    reg [32-1: 0] mem231;
    reg [32-1: 0] mem232;
    reg [32-1: 0] mem233;
    reg [32-1: 0] mem234;
    reg [32-1: 0] mem235;
    reg [32-1: 0] mem236;
    reg [32-1: 0] mem237;
    reg [32-1: 0] mem238;
    reg [32-1: 0] mem239;
    reg [32-1: 0] mem240;
    reg [32-1: 0] mem241;
    reg [32-1: 0] mem242;
    reg [32-1: 0] mem243;
    reg [32-1: 0] mem244;
    reg [32-1: 0] mem245;
    reg [32-1: 0] mem246;
    reg [32-1: 0] mem247;
    reg [32-1: 0] mem248;
    reg [32-1: 0] mem249;
    reg [32-1: 0] mem250;
    reg [32-1: 0] mem251;
    reg [32-1: 0] mem252;
    reg [32-1: 0] mem253;
    reg [32-1: 0] mem254;
    reg [32-1: 0] mem255;
reg [32-1: 0] mem0_n;
    reg [32-1: 0] mem1_n;
    reg [32-1: 0] mem2_n;
    reg [32-1: 0] mem3_n;
    reg [32-1: 0] mem4_n;
    reg [32-1: 0] mem5_n;
    reg [32-1: 0] mem6_n;
    reg [32-1: 0] mem7_n;
    reg [32-1: 0] mem8_n;
    reg [32-1: 0] mem9_n;
    reg [32-1: 0] mem10_n;
    reg [32-1: 0] mem11_n;
    reg [32-1: 0] mem12_n;
    reg [32-1: 0] mem13_n;
    reg [32-1: 0] mem14_n;
    reg [32-1: 0] mem15_n;
    reg [32-1: 0] mem16_n;
    reg [32-1: 0] mem17_n;
    reg [32-1: 0] mem18_n;
    reg [32-1: 0] mem19_n;
    reg [32-1: 0] mem20_n;
    reg [32-1: 0] mem21_n;
    reg [32-1: 0] mem22_n;
    reg [32-1: 0] mem23_n;
    reg [32-1: 0] mem24_n;
    reg [32-1: 0] mem25_n;
    reg [32-1: 0] mem26_n;
    reg [32-1: 0] mem27_n;
    reg [32-1: 0] mem28_n;
    reg [32-1: 0] mem29_n;
    reg [32-1: 0] mem30_n;
    reg [32-1: 0] mem31_n;
    reg [32-1: 0] mem32_n;
    reg [32-1: 0] mem33_n;
    reg [32-1: 0] mem34_n;
    reg [32-1: 0] mem35_n;
    reg [32-1: 0] mem36_n;
    reg [32-1: 0] mem37_n;
    reg [32-1: 0] mem38_n;
    reg [32-1: 0] mem39_n;
    reg [32-1: 0] mem40_n;
    reg [32-1: 0] mem41_n;
    reg [32-1: 0] mem42_n;
    reg [32-1: 0] mem43_n;
    reg [32-1: 0] mem44_n;
    reg [32-1: 0] mem45_n;
    reg [32-1: 0] mem46_n;
    reg [32-1: 0] mem47_n;
    reg [32-1: 0] mem48_n;
    reg [32-1: 0] mem49_n;
    reg [32-1: 0] mem50_n;
    reg [32-1: 0] mem51_n;
    reg [32-1: 0] mem52_n;
    reg [32-1: 0] mem53_n;
    reg [32-1: 0] mem54_n;
    reg [32-1: 0] mem55_n;
    reg [32-1: 0] mem56_n;
    reg [32-1: 0] mem57_n;
    reg [32-1: 0] mem58_n;
    reg [32-1: 0] mem59_n;
    reg [32-1: 0] mem60_n;
    reg [32-1: 0] mem61_n;
    reg [32-1: 0] mem62_n;
    reg [32-1: 0] mem63_n;
    reg [32-1: 0] mem64_n;
    reg [32-1: 0] mem65_n;
    reg [32-1: 0] mem66_n;
    reg [32-1: 0] mem67_n;
    reg [32-1: 0] mem68_n;
    reg [32-1: 0] mem69_n;
    reg [32-1: 0] mem70_n;
    reg [32-1: 0] mem71_n;
    reg [32-1: 0] mem72_n;
    reg [32-1: 0] mem73_n;
    reg [32-1: 0] mem74_n;
    reg [32-1: 0] mem75_n;
    reg [32-1: 0] mem76_n;
    reg [32-1: 0] mem77_n;
    reg [32-1: 0] mem78_n;
    reg [32-1: 0] mem79_n;
    reg [32-1: 0] mem80_n;
    reg [32-1: 0] mem81_n;
    reg [32-1: 0] mem82_n;
    reg [32-1: 0] mem83_n;
    reg [32-1: 0] mem84_n;
    reg [32-1: 0] mem85_n;
    reg [32-1: 0] mem86_n;
    reg [32-1: 0] mem87_n;
    reg [32-1: 0] mem88_n;
    reg [32-1: 0] mem89_n;
    reg [32-1: 0] mem90_n;
    reg [32-1: 0] mem91_n;
    reg [32-1: 0] mem92_n;
    reg [32-1: 0] mem93_n;
    reg [32-1: 0] mem94_n;
    reg [32-1: 0] mem95_n;
    reg [32-1: 0] mem96_n;
    reg [32-1: 0] mem97_n;
    reg [32-1: 0] mem98_n;
    reg [32-1: 0] mem99_n;
    reg [32-1: 0] mem100_n;
    reg [32-1: 0] mem101_n;
    reg [32-1: 0] mem102_n;
    reg [32-1: 0] mem103_n;
    reg [32-1: 0] mem104_n;
    reg [32-1: 0] mem105_n;
    reg [32-1: 0] mem106_n;
    reg [32-1: 0] mem107_n;
    reg [32-1: 0] mem108_n;
    reg [32-1: 0] mem109_n;
    reg [32-1: 0] mem110_n;
    reg [32-1: 0] mem111_n;
    reg [32-1: 0] mem112_n;
    reg [32-1: 0] mem113_n;
    reg [32-1: 0] mem114_n;
    reg [32-1: 0] mem115_n;
    reg [32-1: 0] mem116_n;
    reg [32-1: 0] mem117_n;
    reg [32-1: 0] mem118_n;
    reg [32-1: 0] mem119_n;
    reg [32-1: 0] mem120_n;
    reg [32-1: 0] mem121_n;
    reg [32-1: 0] mem122_n;
    reg [32-1: 0] mem123_n;
    reg [32-1: 0] mem124_n;
    reg [32-1: 0] mem125_n;
    reg [32-1: 0] mem126_n;
    reg [32-1: 0] mem127_n;
    reg [32-1: 0] mem128_n;
    reg [32-1: 0] mem129_n;
    reg [32-1: 0] mem130_n;
    reg [32-1: 0] mem131_n;
    reg [32-1: 0] mem132_n;
    reg [32-1: 0] mem133_n;
    reg [32-1: 0] mem134_n;
    reg [32-1: 0] mem135_n;
    reg [32-1: 0] mem136_n;
    reg [32-1: 0] mem137_n;
    reg [32-1: 0] mem138_n;
    reg [32-1: 0] mem139_n;
    reg [32-1: 0] mem140_n;
    reg [32-1: 0] mem141_n;
    reg [32-1: 0] mem142_n;
    reg [32-1: 0] mem143_n;
    reg [32-1: 0] mem144_n;
    reg [32-1: 0] mem145_n;
    reg [32-1: 0] mem146_n;
    reg [32-1: 0] mem147_n;
    reg [32-1: 0] mem148_n;
    reg [32-1: 0] mem149_n;
    reg [32-1: 0] mem150_n;
    reg [32-1: 0] mem151_n;
    reg [32-1: 0] mem152_n;
    reg [32-1: 0] mem153_n;
    reg [32-1: 0] mem154_n;
    reg [32-1: 0] mem155_n;
    reg [32-1: 0] mem156_n;
    reg [32-1: 0] mem157_n;
    reg [32-1: 0] mem158_n;
    reg [32-1: 0] mem159_n;
    reg [32-1: 0] mem160_n;
    reg [32-1: 0] mem161_n;
    reg [32-1: 0] mem162_n;
    reg [32-1: 0] mem163_n;
    reg [32-1: 0] mem164_n;
    reg [32-1: 0] mem165_n;
    reg [32-1: 0] mem166_n;
    reg [32-1: 0] mem167_n;
    reg [32-1: 0] mem168_n;
    reg [32-1: 0] mem169_n;
    reg [32-1: 0] mem170_n;
    reg [32-1: 0] mem171_n;
    reg [32-1: 0] mem172_n;
    reg [32-1: 0] mem173_n;
    reg [32-1: 0] mem174_n;
    reg [32-1: 0] mem175_n;
    reg [32-1: 0] mem176_n;
    reg [32-1: 0] mem177_n;
    reg [32-1: 0] mem178_n;
    reg [32-1: 0] mem179_n;
    reg [32-1: 0] mem180_n;
    reg [32-1: 0] mem181_n;
    reg [32-1: 0] mem182_n;
    reg [32-1: 0] mem183_n;
    reg [32-1: 0] mem184_n;
    reg [32-1: 0] mem185_n;
    reg [32-1: 0] mem186_n;
    reg [32-1: 0] mem187_n;
    reg [32-1: 0] mem188_n;
    reg [32-1: 0] mem189_n;
    reg [32-1: 0] mem190_n;
    reg [32-1: 0] mem191_n;
    reg [32-1: 0] mem192_n;
    reg [32-1: 0] mem193_n;
    reg [32-1: 0] mem194_n;
    reg [32-1: 0] mem195_n;
    reg [32-1: 0] mem196_n;
    reg [32-1: 0] mem197_n;
    reg [32-1: 0] mem198_n;
    reg [32-1: 0] mem199_n;
    reg [32-1: 0] mem200_n;
    reg [32-1: 0] mem201_n;
    reg [32-1: 0] mem202_n;
    reg [32-1: 0] mem203_n;
    reg [32-1: 0] mem204_n;
    reg [32-1: 0] mem205_n;
    reg [32-1: 0] mem206_n;
    reg [32-1: 0] mem207_n;
    reg [32-1: 0] mem208_n;
    reg [32-1: 0] mem209_n;
    reg [32-1: 0] mem210_n;
    reg [32-1: 0] mem211_n;
    reg [32-1: 0] mem212_n;
    reg [32-1: 0] mem213_n;
    reg [32-1: 0] mem214_n;
    reg [32-1: 0] mem215_n;
    reg [32-1: 0] mem216_n;
    reg [32-1: 0] mem217_n;
    reg [32-1: 0] mem218_n;
    reg [32-1: 0] mem219_n;
    reg [32-1: 0] mem220_n;
    reg [32-1: 0] mem221_n;
    reg [32-1: 0] mem222_n;
    reg [32-1: 0] mem223_n;
    reg [32-1: 0] mem224_n;
    reg [32-1: 0] mem225_n;
    reg [32-1: 0] mem226_n;
    reg [32-1: 0] mem227_n;
    reg [32-1: 0] mem228_n;
    reg [32-1: 0] mem229_n;
    reg [32-1: 0] mem230_n;
    reg [32-1: 0] mem231_n;
    reg [32-1: 0] mem232_n;
    reg [32-1: 0] mem233_n;
    reg [32-1: 0] mem234_n;
    reg [32-1: 0] mem235_n;
    reg [32-1: 0] mem236_n;
    reg [32-1: 0] mem237_n;
    reg [32-1: 0] mem238_n;
    reg [32-1: 0] mem239_n;
    reg [32-1: 0] mem240_n;
    reg [32-1: 0] mem241_n;
    reg [32-1: 0] mem242_n;
    reg [32-1: 0] mem243_n;
    reg [32-1: 0] mem244_n;
    reg [32-1: 0] mem245_n;
    reg [32-1: 0] mem246_n;
    reg [32-1: 0] mem247_n;
    reg [32-1: 0] mem248_n;
    reg [32-1: 0] mem249_n;
    reg [32-1: 0] mem250_n;
    reg [32-1: 0] mem251_n;
    reg [32-1: 0] mem252_n;
    reg [32-1: 0] mem253_n;
    reg [32-1: 0] mem254_n;
    reg [32-1: 0] mem255_n;

always @ (posedge clk) 
    if (~rst_n) begin
        mem0 <= 0;
            mem1 <= 0;
            mem2 <= 0;
            mem3 <= 0;
            mem4 <= 0;
            mem5 <= 0;
            mem6 <= 0;
            mem7 <= 0;
            mem8 <= 0;
            mem9 <= 0;
            mem10 <= 0;
            mem11 <= 0;
            mem12 <= 0;
            mem13 <= 0;
            mem14 <= 0;
            mem15 <= 0;
            mem16 <= 0;
            mem17 <= 0;
            mem18 <= 0;
            mem19 <= 0;
            mem20 <= 0;
            mem21 <= 0;
            mem22 <= 0;
            mem23 <= 0;
            mem24 <= 0;
            mem25 <= 0;
            mem26 <= 0;
            mem27 <= 0;
            mem28 <= 0;
            mem29 <= 0;
            mem30 <= 0;
            mem31 <= 0;
            mem32 <= 0;
            mem33 <= 0;
            mem34 <= 0;
            mem35 <= 0;
            mem36 <= 0;
            mem37 <= 0;
            mem38 <= 0;
            mem39 <= 0;
            mem40 <= 0;
            mem41 <= 0;
            mem42 <= 0;
            mem43 <= 0;
            mem44 <= 0;
            mem45 <= 0;
            mem46 <= 0;
            mem47 <= 0;
            mem48 <= 0;
            mem49 <= 0;
            mem50 <= 0;
            mem51 <= 0;
            mem52 <= 0;
            mem53 <= 0;
            mem54 <= 0;
            mem55 <= 0;
            mem56 <= 0;
            mem57 <= 0;
            mem58 <= 0;
            mem59 <= 0;
            mem60 <= 0;
            mem61 <= 0;
            mem62 <= 0;
            mem63 <= 0;
            mem64 <= 0;
            mem65 <= 0;
            mem66 <= 0;
            mem67 <= 0;
            mem68 <= 0;
            mem69 <= 0;
            mem70 <= 0;
            mem71 <= 0;
            mem72 <= 0;
            mem73 <= 0;
            mem74 <= 0;
            mem75 <= 0;
            mem76 <= 0;
            mem77 <= 0;
            mem78 <= 0;
            mem79 <= 0;
            mem80 <= 0;
            mem81 <= 0;
            mem82 <= 0;
            mem83 <= 0;
            mem84 <= 0;
            mem85 <= 0;
            mem86 <= 0;
            mem87 <= 0;
            mem88 <= 0;
            mem89 <= 0;
            mem90 <= 0;
            mem91 <= 0;
            mem92 <= 0;
            mem93 <= 0;
            mem94 <= 0;
            mem95 <= 0;
            mem96 <= 0;
            mem97 <= 0;
            mem98 <= 0;
            mem99 <= 0;
            mem100 <= 0;
            mem101 <= 0;
            mem102 <= 0;
            mem103 <= 0;
            mem104 <= 0;
            mem105 <= 0;
            mem106 <= 0;
            mem107 <= 0;
            mem108 <= 0;
            mem109 <= 0;
            mem110 <= 0;
            mem111 <= 0;
            mem112 <= 0;
            mem113 <= 0;
            mem114 <= 0;
            mem115 <= 0;
            mem116 <= 0;
            mem117 <= 0;
            mem118 <= 0;
            mem119 <= 0;
            mem120 <= 0;
            mem121 <= 0;
            mem122 <= 0;
            mem123 <= 0;
            mem124 <= 0;
            mem125 <= 0;
            mem126 <= 0;
            mem127 <= 0;
            mem128 <= 0;
            mem129 <= 0;
            mem130 <= 0;
            mem131 <= 0;
            mem132 <= 0;
            mem133 <= 0;
            mem134 <= 0;
            mem135 <= 0;
            mem136 <= 0;
            mem137 <= 0;
            mem138 <= 0;
            mem139 <= 0;
            mem140 <= 0;
            mem141 <= 0;
            mem142 <= 0;
            mem143 <= 0;
            mem144 <= 0;
            mem145 <= 0;
            mem146 <= 0;
            mem147 <= 0;
            mem148 <= 0;
            mem149 <= 0;
            mem150 <= 0;
            mem151 <= 0;
            mem152 <= 0;
            mem153 <= 0;
            mem154 <= 0;
            mem155 <= 0;
            mem156 <= 0;
            mem157 <= 0;
            mem158 <= 0;
            mem159 <= 0;
            mem160 <= 0;
            mem161 <= 0;
            mem162 <= 0;
            mem163 <= 0;
            mem164 <= 0;
            mem165 <= 0;
            mem166 <= 0;
            mem167 <= 0;
            mem168 <= 0;
            mem169 <= 0;
            mem170 <= 0;
            mem171 <= 0;
            mem172 <= 0;
            mem173 <= 0;
            mem174 <= 0;
            mem175 <= 0;
            mem176 <= 0;
            mem177 <= 0;
            mem178 <= 0;
            mem179 <= 0;
            mem180 <= 0;
            mem181 <= 0;
            mem182 <= 0;
            mem183 <= 0;
            mem184 <= 0;
            mem185 <= 0;
            mem186 <= 0;
            mem187 <= 0;
            mem188 <= 0;
            mem189 <= 0;
            mem190 <= 0;
            mem191 <= 0;
            mem192 <= 0;
            mem193 <= 0;
            mem194 <= 0;
            mem195 <= 0;
            mem196 <= 0;
            mem197 <= 0;
            mem198 <= 0;
            mem199 <= 0;
            mem200 <= 0;
            mem201 <= 0;
            mem202 <= 0;
            mem203 <= 0;
            mem204 <= 0;
            mem205 <= 0;
            mem206 <= 0;
            mem207 <= 0;
            mem208 <= 0;
            mem209 <= 0;
            mem210 <= 0;
            mem211 <= 0;
            mem212 <= 0;
            mem213 <= 0;
            mem214 <= 0;
            mem215 <= 0;
            mem216 <= 0;
            mem217 <= 0;
            mem218 <= 0;
            mem219 <= 0;
            mem220 <= 0;
            mem221 <= 0;
            mem222 <= 0;
            mem223 <= 0;
            mem224 <= 0;
            mem225 <= 0;
            mem226 <= 0;
            mem227 <= 0;
            mem228 <= 0;
            mem229 <= 0;
            mem230 <= 0;
            mem231 <= 0;
            mem232 <= 0;
            mem233 <= 0;
            mem234 <= 0;
            mem235 <= 0;
            mem236 <= 0;
            mem237 <= 0;
            mem238 <= 0;
            mem239 <= 0;
            mem240 <= 0;
            mem241 <= 0;
            mem242 <= 0;
            mem243 <= 0;
            mem244 <= 0;
            mem245 <= 0;
            mem246 <= 0;
            mem247 <= 0;
            mem248 <= 0;
            mem249 <= 0;
            mem250 <= 0;
            mem251 <= 0;
            mem252 <= 0;
            mem253 <= 0;
            mem254 <= 0;
            mem255 <= 0;
    end
    else begin

        mem0 <= mem0_n;
            mem1 <= mem1_n;
            mem2 <= mem2_n;
            mem3 <= mem3_n;
            mem4 <= mem4_n;
            mem5 <= mem5_n;
            mem6 <= mem6_n;
            mem7 <= mem7_n;
            mem8 <= mem8_n;
            mem9 <= mem9_n;
            mem10 <= mem10_n;
            mem11 <= mem11_n;
            mem12 <= mem12_n;
            mem13 <= mem13_n;
            mem14 <= mem14_n;
            mem15 <= mem15_n;
            mem16 <= mem16_n;
            mem17 <= mem17_n;
            mem18 <= mem18_n;
            mem19 <= mem19_n;
            mem20 <= mem20_n;
            mem21 <= mem21_n;
            mem22 <= mem22_n;
            mem23 <= mem23_n;
            mem24 <= mem24_n;
            mem25 <= mem25_n;
            mem26 <= mem26_n;
            mem27 <= mem27_n;
            mem28 <= mem28_n;
            mem29 <= mem29_n;
            mem30 <= mem30_n;
            mem31 <= mem31_n;
            mem32 <= mem32_n;
            mem33 <= mem33_n;
            mem34 <= mem34_n;
            mem35 <= mem35_n;
            mem36 <= mem36_n;
            mem37 <= mem37_n;
            mem38 <= mem38_n;
            mem39 <= mem39_n;
            mem40 <= mem40_n;
            mem41 <= mem41_n;
            mem42 <= mem42_n;
            mem43 <= mem43_n;
            mem44 <= mem44_n;
            mem45 <= mem45_n;
            mem46 <= mem46_n;
            mem47 <= mem47_n;
            mem48 <= mem48_n;
            mem49 <= mem49_n;
            mem50 <= mem50_n;
            mem51 <= mem51_n;
            mem52 <= mem52_n;
            mem53 <= mem53_n;
            mem54 <= mem54_n;
            mem55 <= mem55_n;
            mem56 <= mem56_n;
            mem57 <= mem57_n;
            mem58 <= mem58_n;
            mem59 <= mem59_n;
            mem60 <= mem60_n;
            mem61 <= mem61_n;
            mem62 <= mem62_n;
            mem63 <= mem63_n;
            mem64 <= mem64_n;
            mem65 <= mem65_n;
            mem66 <= mem66_n;
            mem67 <= mem67_n;
            mem68 <= mem68_n;
            mem69 <= mem69_n;
            mem70 <= mem70_n;
            mem71 <= mem71_n;
            mem72 <= mem72_n;
            mem73 <= mem73_n;
            mem74 <= mem74_n;
            mem75 <= mem75_n;
            mem76 <= mem76_n;
            mem77 <= mem77_n;
            mem78 <= mem78_n;
            mem79 <= mem79_n;
            mem80 <= mem80_n;
            mem81 <= mem81_n;
            mem82 <= mem82_n;
            mem83 <= mem83_n;
            mem84 <= mem84_n;
            mem85 <= mem85_n;
            mem86 <= mem86_n;
            mem87 <= mem87_n;
            mem88 <= mem88_n;
            mem89 <= mem89_n;
            mem90 <= mem90_n;
            mem91 <= mem91_n;
            mem92 <= mem92_n;
            mem93 <= mem93_n;
            mem94 <= mem94_n;
            mem95 <= mem95_n;
            mem96 <= mem96_n;
            mem97 <= mem97_n;
            mem98 <= mem98_n;
            mem99 <= mem99_n;
            mem100 <= mem100_n;
            mem101 <= mem101_n;
            mem102 <= mem102_n;
            mem103 <= mem103_n;
            mem104 <= mem104_n;
            mem105 <= mem105_n;
            mem106 <= mem106_n;
            mem107 <= mem107_n;
            mem108 <= mem108_n;
            mem109 <= mem109_n;
            mem110 <= mem110_n;
            mem111 <= mem111_n;
            mem112 <= mem112_n;
            mem113 <= mem113_n;
            mem114 <= mem114_n;
            mem115 <= mem115_n;
            mem116 <= mem116_n;
            mem117 <= mem117_n;
            mem118 <= mem118_n;
            mem119 <= mem119_n;
            mem120 <= mem120_n;
            mem121 <= mem121_n;
            mem122 <= mem122_n;
            mem123 <= mem123_n;
            mem124 <= mem124_n;
            mem125 <= mem125_n;
            mem126 <= mem126_n;
            mem127 <= mem127_n;
            mem128 <= mem128_n;
            mem129 <= mem129_n;
            mem130 <= mem130_n;
            mem131 <= mem131_n;
            mem132 <= mem132_n;
            mem133 <= mem133_n;
            mem134 <= mem134_n;
            mem135 <= mem135_n;
            mem136 <= mem136_n;
            mem137 <= mem137_n;
            mem138 <= mem138_n;
            mem139 <= mem139_n;
            mem140 <= mem140_n;
            mem141 <= mem141_n;
            mem142 <= mem142_n;
            mem143 <= mem143_n;
            mem144 <= mem144_n;
            mem145 <= mem145_n;
            mem146 <= mem146_n;
            mem147 <= mem147_n;
            mem148 <= mem148_n;
            mem149 <= mem149_n;
            mem150 <= mem150_n;
            mem151 <= mem151_n;
            mem152 <= mem152_n;
            mem153 <= mem153_n;
            mem154 <= mem154_n;
            mem155 <= mem155_n;
            mem156 <= mem156_n;
            mem157 <= mem157_n;
            mem158 <= mem158_n;
            mem159 <= mem159_n;
            mem160 <= mem160_n;
            mem161 <= mem161_n;
            mem162 <= mem162_n;
            mem163 <= mem163_n;
            mem164 <= mem164_n;
            mem165 <= mem165_n;
            mem166 <= mem166_n;
            mem167 <= mem167_n;
            mem168 <= mem168_n;
            mem169 <= mem169_n;
            mem170 <= mem170_n;
            mem171 <= mem171_n;
            mem172 <= mem172_n;
            mem173 <= mem173_n;
            mem174 <= mem174_n;
            mem175 <= mem175_n;
            mem176 <= mem176_n;
            mem177 <= mem177_n;
            mem178 <= mem178_n;
            mem179 <= mem179_n;
            mem180 <= mem180_n;
            mem181 <= mem181_n;
            mem182 <= mem182_n;
            mem183 <= mem183_n;
            mem184 <= mem184_n;
            mem185 <= mem185_n;
            mem186 <= mem186_n;
            mem187 <= mem187_n;
            mem188 <= mem188_n;
            mem189 <= mem189_n;
            mem190 <= mem190_n;
            mem191 <= mem191_n;
            mem192 <= mem192_n;
            mem193 <= mem193_n;
            mem194 <= mem194_n;
            mem195 <= mem195_n;
            mem196 <= mem196_n;
            mem197 <= mem197_n;
            mem198 <= mem198_n;
            mem199 <= mem199_n;
            mem200 <= mem200_n;
            mem201 <= mem201_n;
            mem202 <= mem202_n;
            mem203 <= mem203_n;
            mem204 <= mem204_n;
            mem205 <= mem205_n;
            mem206 <= mem206_n;
            mem207 <= mem207_n;
            mem208 <= mem208_n;
            mem209 <= mem209_n;
            mem210 <= mem210_n;
            mem211 <= mem211_n;
            mem212 <= mem212_n;
            mem213 <= mem213_n;
            mem214 <= mem214_n;
            mem215 <= mem215_n;
            mem216 <= mem216_n;
            mem217 <= mem217_n;
            mem218 <= mem218_n;
            mem219 <= mem219_n;
            mem220 <= mem220_n;
            mem221 <= mem221_n;
            mem222 <= mem222_n;
            mem223 <= mem223_n;
            mem224 <= mem224_n;
            mem225 <= mem225_n;
            mem226 <= mem226_n;
            mem227 <= mem227_n;
            mem228 <= mem228_n;
            mem229 <= mem229_n;
            mem230 <= mem230_n;
            mem231 <= mem231_n;
            mem232 <= mem232_n;
            mem233 <= mem233_n;
            mem234 <= mem234_n;
            mem235 <= mem235_n;
            mem236 <= mem236_n;
            mem237 <= mem237_n;
            mem238 <= mem238_n;
            mem239 <= mem239_n;
            mem240 <= mem240_n;
            mem241 <= mem241_n;
            mem242 <= mem242_n;
            mem243 <= mem243_n;
            mem244 <= mem244_n;
            mem245 <= mem245_n;
            mem246 <= mem246_n;
            mem247 <= mem247_n;
            mem248 <= mem248_n;
            mem249 <= mem249_n;
            mem250 <= mem250_n;
            mem251 <= mem251_n;
            mem252 <= mem252_n;
            mem253 <= mem253_n;
            mem254 <= mem254_n;
            mem255 <= mem255_n;
    end

always@* begin
    rdata = 0;
    case (addr)

        0: rdata = mem0;
            1: rdata = mem1;
            2: rdata = mem2;
            3: rdata = mem3;
            4: rdata = mem4;
            5: rdata = mem5;
            6: rdata = mem6;
            7: rdata = mem7;
            8: rdata = mem8;
            9: rdata = mem9;
            10: rdata = mem10;
            11: rdata = mem11;
            12: rdata = mem12;
            13: rdata = mem13;
            14: rdata = mem14;
            15: rdata = mem15;
            16: rdata = mem16;
            17: rdata = mem17;
            18: rdata = mem18;
            19: rdata = mem19;
            20: rdata = mem20;
            21: rdata = mem21;
            22: rdata = mem22;
            23: rdata = mem23;
            24: rdata = mem24;
            25: rdata = mem25;
            26: rdata = mem26;
            27: rdata = mem27;
            28: rdata = mem28;
            29: rdata = mem29;
            30: rdata = mem30;
            31: rdata = mem31;
            32: rdata = mem32;
            33: rdata = mem33;
            34: rdata = mem34;
            35: rdata = mem35;
            36: rdata = mem36;
            37: rdata = mem37;
            38: rdata = mem38;
            39: rdata = mem39;
            40: rdata = mem40;
            41: rdata = mem41;
            42: rdata = mem42;
            43: rdata = mem43;
            44: rdata = mem44;
            45: rdata = mem45;
            46: rdata = mem46;
            47: rdata = mem47;
            48: rdata = mem48;
            49: rdata = mem49;
            50: rdata = mem50;
            51: rdata = mem51;
            52: rdata = mem52;
            53: rdata = mem53;
            54: rdata = mem54;
            55: rdata = mem55;
            56: rdata = mem56;
            57: rdata = mem57;
            58: rdata = mem58;
            59: rdata = mem59;
            60: rdata = mem60;
            61: rdata = mem61;
            62: rdata = mem62;
            63: rdata = mem63;
            64: rdata = mem64;
            65: rdata = mem65;
            66: rdata = mem66;
            67: rdata = mem67;
            68: rdata = mem68;
            69: rdata = mem69;
            70: rdata = mem70;
            71: rdata = mem71;
            72: rdata = mem72;
            73: rdata = mem73;
            74: rdata = mem74;
            75: rdata = mem75;
            76: rdata = mem76;
            77: rdata = mem77;
            78: rdata = mem78;
            79: rdata = mem79;
            80: rdata = mem80;
            81: rdata = mem81;
            82: rdata = mem82;
            83: rdata = mem83;
            84: rdata = mem84;
            85: rdata = mem85;
            86: rdata = mem86;
            87: rdata = mem87;
            88: rdata = mem88;
            89: rdata = mem89;
            90: rdata = mem90;
            91: rdata = mem91;
            92: rdata = mem92;
            93: rdata = mem93;
            94: rdata = mem94;
            95: rdata = mem95;
            96: rdata = mem96;
            97: rdata = mem97;
            98: rdata = mem98;
            99: rdata = mem99;
            100: rdata = mem100;
            101: rdata = mem101;
            102: rdata = mem102;
            103: rdata = mem103;
            104: rdata = mem104;
            105: rdata = mem105;
            106: rdata = mem106;
            107: rdata = mem107;
            108: rdata = mem108;
            109: rdata = mem109;
            110: rdata = mem110;
            111: rdata = mem111;
            112: rdata = mem112;
            113: rdata = mem113;
            114: rdata = mem114;
            115: rdata = mem115;
            116: rdata = mem116;
            117: rdata = mem117;
            118: rdata = mem118;
            119: rdata = mem119;
            120: rdata = mem120;
            121: rdata = mem121;
            122: rdata = mem122;
            123: rdata = mem123;
            124: rdata = mem124;
            125: rdata = mem125;
            126: rdata = mem126;
            127: rdata = mem127;
            128: rdata = mem128;
            129: rdata = mem129;
            130: rdata = mem130;
            131: rdata = mem131;
            132: rdata = mem132;
            133: rdata = mem133;
            134: rdata = mem134;
            135: rdata = mem135;
            136: rdata = mem136;
            137: rdata = mem137;
            138: rdata = mem138;
            139: rdata = mem139;
            140: rdata = mem140;
            141: rdata = mem141;
            142: rdata = mem142;
            143: rdata = mem143;
            144: rdata = mem144;
            145: rdata = mem145;
            146: rdata = mem146;
            147: rdata = mem147;
            148: rdata = mem148;
            149: rdata = mem149;
            150: rdata = mem150;
            151: rdata = mem151;
            152: rdata = mem152;
            153: rdata = mem153;
            154: rdata = mem154;
            155: rdata = mem155;
            156: rdata = mem156;
            157: rdata = mem157;
            158: rdata = mem158;
            159: rdata = mem159;
            160: rdata = mem160;
            161: rdata = mem161;
            162: rdata = mem162;
            163: rdata = mem163;
            164: rdata = mem164;
            165: rdata = mem165;
            166: rdata = mem166;
            167: rdata = mem167;
            168: rdata = mem168;
            169: rdata = mem169;
            170: rdata = mem170;
            171: rdata = mem171;
            172: rdata = mem172;
            173: rdata = mem173;
            174: rdata = mem174;
            175: rdata = mem175;
            176: rdata = mem176;
            177: rdata = mem177;
            178: rdata = mem178;
            179: rdata = mem179;
            180: rdata = mem180;
            181: rdata = mem181;
            182: rdata = mem182;
            183: rdata = mem183;
            184: rdata = mem184;
            185: rdata = mem185;
            186: rdata = mem186;
            187: rdata = mem187;
            188: rdata = mem188;
            189: rdata = mem189;
            190: rdata = mem190;
            191: rdata = mem191;
            192: rdata = mem192;
            193: rdata = mem193;
            194: rdata = mem194;
            195: rdata = mem195;
            196: rdata = mem196;
            197: rdata = mem197;
            198: rdata = mem198;
            199: rdata = mem199;
            200: rdata = mem200;
            201: rdata = mem201;
            202: rdata = mem202;
            203: rdata = mem203;
            204: rdata = mem204;
            205: rdata = mem205;
            206: rdata = mem206;
            207: rdata = mem207;
            208: rdata = mem208;
            209: rdata = mem209;
            210: rdata = mem210;
            211: rdata = mem211;
            212: rdata = mem212;
            213: rdata = mem213;
            214: rdata = mem214;
            215: rdata = mem215;
            216: rdata = mem216;
            217: rdata = mem217;
            218: rdata = mem218;
            219: rdata = mem219;
            220: rdata = mem220;
            221: rdata = mem221;
            222: rdata = mem222;
            223: rdata = mem223;
            224: rdata = mem224;
            225: rdata = mem225;
            226: rdata = mem226;
            227: rdata = mem227;
            228: rdata = mem228;
            229: rdata = mem229;
            230: rdata = mem230;
            231: rdata = mem231;
            232: rdata = mem232;
            233: rdata = mem233;
            234: rdata = mem234;
            235: rdata = mem235;
            236: rdata = mem236;
            237: rdata = mem237;
            238: rdata = mem238;
            239: rdata = mem239;
            240: rdata = mem240;
            241: rdata = mem241;
            242: rdata = mem242;
            243: rdata = mem243;
            244: rdata = mem244;
            245: rdata = mem245;
            246: rdata = mem246;
            247: rdata = mem247;
            248: rdata = mem248;
            249: rdata = mem249;
            250: rdata = mem250;
            251: rdata = mem251;
            252: rdata = mem252;
            253: rdata = mem253;
            254: rdata = mem254;
            255: rdata = mem255;
    endcase
end

always @(*) begin

        mem0_n = (wen && ( 0 == addr))? wdata : mem0; 
            mem1_n = (wen && ( 1 == addr))? wdata : mem1; 
            mem2_n = (wen && ( 2 == addr))? wdata : mem2; 
            mem3_n = (wen && ( 3 == addr))? wdata : mem3; 
            mem4_n = (wen && ( 4 == addr))? wdata : mem4; 
            mem5_n = (wen && ( 5 == addr))? wdata : mem5; 
            mem6_n = (wen && ( 6 == addr))? wdata : mem6; 
            mem7_n = (wen && ( 7 == addr))? wdata : mem7; 
            mem8_n = (wen && ( 8 == addr))? wdata : mem8; 
            mem9_n = (wen && ( 9 == addr))? wdata : mem9; 
            mem10_n = (wen && ( 10 == addr))? wdata : mem10; 
            mem11_n = (wen && ( 11 == addr))? wdata : mem11; 
            mem12_n = (wen && ( 12 == addr))? wdata : mem12; 
            mem13_n = (wen && ( 13 == addr))? wdata : mem13; 
            mem14_n = (wen && ( 14 == addr))? wdata : mem14; 
            mem15_n = (wen && ( 15 == addr))? wdata : mem15; 
            mem16_n = (wen && ( 16 == addr))? wdata : mem16; 
            mem17_n = (wen && ( 17 == addr))? wdata : mem17; 
            mem18_n = (wen && ( 18 == addr))? wdata : mem18; 
            mem19_n = (wen && ( 19 == addr))? wdata : mem19; 
            mem20_n = (wen && ( 20 == addr))? wdata : mem20; 
            mem21_n = (wen && ( 21 == addr))? wdata : mem21; 
            mem22_n = (wen && ( 22 == addr))? wdata : mem22; 
            mem23_n = (wen && ( 23 == addr))? wdata : mem23; 
            mem24_n = (wen && ( 24 == addr))? wdata : mem24; 
            mem25_n = (wen && ( 25 == addr))? wdata : mem25; 
            mem26_n = (wen && ( 26 == addr))? wdata : mem26; 
            mem27_n = (wen && ( 27 == addr))? wdata : mem27; 
            mem28_n = (wen && ( 28 == addr))? wdata : mem28; 
            mem29_n = (wen && ( 29 == addr))? wdata : mem29; 
            mem30_n = (wen && ( 30 == addr))? wdata : mem30; 
            mem31_n = (wen && ( 31 == addr))? wdata : mem31; 
            mem32_n = (wen && ( 32 == addr))? wdata : mem32; 
            mem33_n = (wen && ( 33 == addr))? wdata : mem33; 
            mem34_n = (wen && ( 34 == addr))? wdata : mem34; 
            mem35_n = (wen && ( 35 == addr))? wdata : mem35; 
            mem36_n = (wen && ( 36 == addr))? wdata : mem36; 
            mem37_n = (wen && ( 37 == addr))? wdata : mem37; 
            mem38_n = (wen && ( 38 == addr))? wdata : mem38; 
            mem39_n = (wen && ( 39 == addr))? wdata : mem39; 
            mem40_n = (wen && ( 40 == addr))? wdata : mem40; 
            mem41_n = (wen && ( 41 == addr))? wdata : mem41; 
            mem42_n = (wen && ( 42 == addr))? wdata : mem42; 
            mem43_n = (wen && ( 43 == addr))? wdata : mem43; 
            mem44_n = (wen && ( 44 == addr))? wdata : mem44; 
            mem45_n = (wen && ( 45 == addr))? wdata : mem45; 
            mem46_n = (wen && ( 46 == addr))? wdata : mem46; 
            mem47_n = (wen && ( 47 == addr))? wdata : mem47; 
            mem48_n = (wen && ( 48 == addr))? wdata : mem48; 
            mem49_n = (wen && ( 49 == addr))? wdata : mem49; 
            mem50_n = (wen && ( 50 == addr))? wdata : mem50; 
            mem51_n = (wen && ( 51 == addr))? wdata : mem51; 
            mem52_n = (wen && ( 52 == addr))? wdata : mem52; 
            mem53_n = (wen && ( 53 == addr))? wdata : mem53; 
            mem54_n = (wen && ( 54 == addr))? wdata : mem54; 
            mem55_n = (wen && ( 55 == addr))? wdata : mem55; 
            mem56_n = (wen && ( 56 == addr))? wdata : mem56; 
            mem57_n = (wen && ( 57 == addr))? wdata : mem57; 
            mem58_n = (wen && ( 58 == addr))? wdata : mem58; 
            mem59_n = (wen && ( 59 == addr))? wdata : mem59; 
            mem60_n = (wen && ( 60 == addr))? wdata : mem60; 
            mem61_n = (wen && ( 61 == addr))? wdata : mem61; 
            mem62_n = (wen && ( 62 == addr))? wdata : mem62; 
            mem63_n = (wen && ( 63 == addr))? wdata : mem63; 
            mem64_n = (wen && ( 64 == addr))? wdata : mem64; 
            mem65_n = (wen && ( 65 == addr))? wdata : mem65; 
            mem66_n = (wen && ( 66 == addr))? wdata : mem66; 
            mem67_n = (wen && ( 67 == addr))? wdata : mem67; 
            mem68_n = (wen && ( 68 == addr))? wdata : mem68; 
            mem69_n = (wen && ( 69 == addr))? wdata : mem69; 
            mem70_n = (wen && ( 70 == addr))? wdata : mem70; 
            mem71_n = (wen && ( 71 == addr))? wdata : mem71; 
            mem72_n = (wen && ( 72 == addr))? wdata : mem72; 
            mem73_n = (wen && ( 73 == addr))? wdata : mem73; 
            mem74_n = (wen && ( 74 == addr))? wdata : mem74; 
            mem75_n = (wen && ( 75 == addr))? wdata : mem75; 
            mem76_n = (wen && ( 76 == addr))? wdata : mem76; 
            mem77_n = (wen && ( 77 == addr))? wdata : mem77; 
            mem78_n = (wen && ( 78 == addr))? wdata : mem78; 
            mem79_n = (wen && ( 79 == addr))? wdata : mem79; 
            mem80_n = (wen && ( 80 == addr))? wdata : mem80; 
            mem81_n = (wen && ( 81 == addr))? wdata : mem81; 
            mem82_n = (wen && ( 82 == addr))? wdata : mem82; 
            mem83_n = (wen && ( 83 == addr))? wdata : mem83; 
            mem84_n = (wen && ( 84 == addr))? wdata : mem84; 
            mem85_n = (wen && ( 85 == addr))? wdata : mem85; 
            mem86_n = (wen && ( 86 == addr))? wdata : mem86; 
            mem87_n = (wen && ( 87 == addr))? wdata : mem87; 
            mem88_n = (wen && ( 88 == addr))? wdata : mem88; 
            mem89_n = (wen && ( 89 == addr))? wdata : mem89; 
            mem90_n = (wen && ( 90 == addr))? wdata : mem90; 
            mem91_n = (wen && ( 91 == addr))? wdata : mem91; 
            mem92_n = (wen && ( 92 == addr))? wdata : mem92; 
            mem93_n = (wen && ( 93 == addr))? wdata : mem93; 
            mem94_n = (wen && ( 94 == addr))? wdata : mem94; 
            mem95_n = (wen && ( 95 == addr))? wdata : mem95; 
            mem96_n = (wen && ( 96 == addr))? wdata : mem96; 
            mem97_n = (wen && ( 97 == addr))? wdata : mem97; 
            mem98_n = (wen && ( 98 == addr))? wdata : mem98; 
            mem99_n = (wen && ( 99 == addr))? wdata : mem99; 
            mem100_n = (wen && ( 100 == addr))? wdata : mem100; 
            mem101_n = (wen && ( 101 == addr))? wdata : mem101; 
            mem102_n = (wen && ( 102 == addr))? wdata : mem102; 
            mem103_n = (wen && ( 103 == addr))? wdata : mem103; 
            mem104_n = (wen && ( 104 == addr))? wdata : mem104; 
            mem105_n = (wen && ( 105 == addr))? wdata : mem105; 
            mem106_n = (wen && ( 106 == addr))? wdata : mem106; 
            mem107_n = (wen && ( 107 == addr))? wdata : mem107; 
            mem108_n = (wen && ( 108 == addr))? wdata : mem108; 
            mem109_n = (wen && ( 109 == addr))? wdata : mem109; 
            mem110_n = (wen && ( 110 == addr))? wdata : mem110; 
            mem111_n = (wen && ( 111 == addr))? wdata : mem111; 
            mem112_n = (wen && ( 112 == addr))? wdata : mem112; 
            mem113_n = (wen && ( 113 == addr))? wdata : mem113; 
            mem114_n = (wen && ( 114 == addr))? wdata : mem114; 
            mem115_n = (wen && ( 115 == addr))? wdata : mem115; 
            mem116_n = (wen && ( 116 == addr))? wdata : mem116; 
            mem117_n = (wen && ( 117 == addr))? wdata : mem117; 
            mem118_n = (wen && ( 118 == addr))? wdata : mem118; 
            mem119_n = (wen && ( 119 == addr))? wdata : mem119; 
            mem120_n = (wen && ( 120 == addr))? wdata : mem120; 
            mem121_n = (wen && ( 121 == addr))? wdata : mem121; 
            mem122_n = (wen && ( 122 == addr))? wdata : mem122; 
            mem123_n = (wen && ( 123 == addr))? wdata : mem123; 
            mem124_n = (wen && ( 124 == addr))? wdata : mem124; 
            mem125_n = (wen && ( 125 == addr))? wdata : mem125; 
            mem126_n = (wen && ( 126 == addr))? wdata : mem126; 
            mem127_n = (wen && ( 127 == addr))? wdata : mem127; 
            mem128_n = (wen && ( 128 == addr))? wdata : mem128; 
            mem129_n = (wen && ( 129 == addr))? wdata : mem129; 
            mem130_n = (wen && ( 130 == addr))? wdata : mem130; 
            mem131_n = (wen && ( 131 == addr))? wdata : mem131; 
            mem132_n = (wen && ( 132 == addr))? wdata : mem132; 
            mem133_n = (wen && ( 133 == addr))? wdata : mem133; 
            mem134_n = (wen && ( 134 == addr))? wdata : mem134; 
            mem135_n = (wen && ( 135 == addr))? wdata : mem135; 
            mem136_n = (wen && ( 136 == addr))? wdata : mem136; 
            mem137_n = (wen && ( 137 == addr))? wdata : mem137; 
            mem138_n = (wen && ( 138 == addr))? wdata : mem138; 
            mem139_n = (wen && ( 139 == addr))? wdata : mem139; 
            mem140_n = (wen && ( 140 == addr))? wdata : mem140; 
            mem141_n = (wen && ( 141 == addr))? wdata : mem141; 
            mem142_n = (wen && ( 142 == addr))? wdata : mem142; 
            mem143_n = (wen && ( 143 == addr))? wdata : mem143; 
            mem144_n = (wen && ( 144 == addr))? wdata : mem144; 
            mem145_n = (wen && ( 145 == addr))? wdata : mem145; 
            mem146_n = (wen && ( 146 == addr))? wdata : mem146; 
            mem147_n = (wen && ( 147 == addr))? wdata : mem147; 
            mem148_n = (wen && ( 148 == addr))? wdata : mem148; 
            mem149_n = (wen && ( 149 == addr))? wdata : mem149; 
            mem150_n = (wen && ( 150 == addr))? wdata : mem150; 
            mem151_n = (wen && ( 151 == addr))? wdata : mem151; 
            mem152_n = (wen && ( 152 == addr))? wdata : mem152; 
            mem153_n = (wen && ( 153 == addr))? wdata : mem153; 
            mem154_n = (wen && ( 154 == addr))? wdata : mem154; 
            mem155_n = (wen && ( 155 == addr))? wdata : mem155; 
            mem156_n = (wen && ( 156 == addr))? wdata : mem156; 
            mem157_n = (wen && ( 157 == addr))? wdata : mem157; 
            mem158_n = (wen && ( 158 == addr))? wdata : mem158; 
            mem159_n = (wen && ( 159 == addr))? wdata : mem159; 
            mem160_n = (wen && ( 160 == addr))? wdata : mem160; 
            mem161_n = (wen && ( 161 == addr))? wdata : mem161; 
            mem162_n = (wen && ( 162 == addr))? wdata : mem162; 
            mem163_n = (wen && ( 163 == addr))? wdata : mem163; 
            mem164_n = (wen && ( 164 == addr))? wdata : mem164; 
            mem165_n = (wen && ( 165 == addr))? wdata : mem165; 
            mem166_n = (wen && ( 166 == addr))? wdata : mem166; 
            mem167_n = (wen && ( 167 == addr))? wdata : mem167; 
            mem168_n = (wen && ( 168 == addr))? wdata : mem168; 
            mem169_n = (wen && ( 169 == addr))? wdata : mem169; 
            mem170_n = (wen && ( 170 == addr))? wdata : mem170; 
            mem171_n = (wen && ( 171 == addr))? wdata : mem171; 
            mem172_n = (wen && ( 172 == addr))? wdata : mem172; 
            mem173_n = (wen && ( 173 == addr))? wdata : mem173; 
            mem174_n = (wen && ( 174 == addr))? wdata : mem174; 
            mem175_n = (wen && ( 175 == addr))? wdata : mem175; 
            mem176_n = (wen && ( 176 == addr))? wdata : mem176; 
            mem177_n = (wen && ( 177 == addr))? wdata : mem177; 
            mem178_n = (wen && ( 178 == addr))? wdata : mem178; 
            mem179_n = (wen && ( 179 == addr))? wdata : mem179; 
            mem180_n = (wen && ( 180 == addr))? wdata : mem180; 
            mem181_n = (wen && ( 181 == addr))? wdata : mem181; 
            mem182_n = (wen && ( 182 == addr))? wdata : mem182; 
            mem183_n = (wen && ( 183 == addr))? wdata : mem183; 
            mem184_n = (wen && ( 184 == addr))? wdata : mem184; 
            mem185_n = (wen && ( 185 == addr))? wdata : mem185; 
            mem186_n = (wen && ( 186 == addr))? wdata : mem186; 
            mem187_n = (wen && ( 187 == addr))? wdata : mem187; 
            mem188_n = (wen && ( 188 == addr))? wdata : mem188; 
            mem189_n = (wen && ( 189 == addr))? wdata : mem189; 
            mem190_n = (wen && ( 190 == addr))? wdata : mem190; 
            mem191_n = (wen && ( 191 == addr))? wdata : mem191; 
            mem192_n = (wen && ( 192 == addr))? wdata : mem192; 
            mem193_n = (wen && ( 193 == addr))? wdata : mem193; 
            mem194_n = (wen && ( 194 == addr))? wdata : mem194; 
            mem195_n = (wen && ( 195 == addr))? wdata : mem195; 
            mem196_n = (wen && ( 196 == addr))? wdata : mem196; 
            mem197_n = (wen && ( 197 == addr))? wdata : mem197; 
            mem198_n = (wen && ( 198 == addr))? wdata : mem198; 
            mem199_n = (wen && ( 199 == addr))? wdata : mem199; 
            mem200_n = (wen && ( 200 == addr))? wdata : mem200; 
            mem201_n = (wen && ( 201 == addr))? wdata : mem201; 
            mem202_n = (wen && ( 202 == addr))? wdata : mem202; 
            mem203_n = (wen && ( 203 == addr))? wdata : mem203; 
            mem204_n = (wen && ( 204 == addr))? wdata : mem204; 
            mem205_n = (wen && ( 205 == addr))? wdata : mem205; 
            mem206_n = (wen && ( 206 == addr))? wdata : mem206; 
            mem207_n = (wen && ( 207 == addr))? wdata : mem207; 
            mem208_n = (wen && ( 208 == addr))? wdata : mem208; 
            mem209_n = (wen && ( 209 == addr))? wdata : mem209; 
            mem210_n = (wen && ( 210 == addr))? wdata : mem210; 
            mem211_n = (wen && ( 211 == addr))? wdata : mem211; 
            mem212_n = (wen && ( 212 == addr))? wdata : mem212; 
            mem213_n = (wen && ( 213 == addr))? wdata : mem213; 
            mem214_n = (wen && ( 214 == addr))? wdata : mem214; 
            mem215_n = (wen && ( 215 == addr))? wdata : mem215; 
            mem216_n = (wen && ( 216 == addr))? wdata : mem216; 
            mem217_n = (wen && ( 217 == addr))? wdata : mem217; 
            mem218_n = (wen && ( 218 == addr))? wdata : mem218; 
            mem219_n = (wen && ( 219 == addr))? wdata : mem219; 
            mem220_n = (wen && ( 220 == addr))? wdata : mem220; 
            mem221_n = (wen && ( 221 == addr))? wdata : mem221; 
            mem222_n = (wen && ( 222 == addr))? wdata : mem222; 
            mem223_n = (wen && ( 223 == addr))? wdata : mem223; 
            mem224_n = (wen && ( 224 == addr))? wdata : mem224; 
            mem225_n = (wen && ( 225 == addr))? wdata : mem225; 
            mem226_n = (wen && ( 226 == addr))? wdata : mem226; 
            mem227_n = (wen && ( 227 == addr))? wdata : mem227; 
            mem228_n = (wen && ( 228 == addr))? wdata : mem228; 
            mem229_n = (wen && ( 229 == addr))? wdata : mem229; 
            mem230_n = (wen && ( 230 == addr))? wdata : mem230; 
            mem231_n = (wen && ( 231 == addr))? wdata : mem231; 
            mem232_n = (wen && ( 232 == addr))? wdata : mem232; 
            mem233_n = (wen && ( 233 == addr))? wdata : mem233; 
            mem234_n = (wen && ( 234 == addr))? wdata : mem234; 
            mem235_n = (wen && ( 235 == addr))? wdata : mem235; 
            mem236_n = (wen && ( 236 == addr))? wdata : mem236; 
            mem237_n = (wen && ( 237 == addr))? wdata : mem237; 
            mem238_n = (wen && ( 238 == addr))? wdata : mem238; 
            mem239_n = (wen && ( 239 == addr))? wdata : mem239; 
            mem240_n = (wen && ( 240 == addr))? wdata : mem240; 
            mem241_n = (wen && ( 241 == addr))? wdata : mem241; 
            mem242_n = (wen && ( 242 == addr))? wdata : mem242; 
            mem243_n = (wen && ( 243 == addr))? wdata : mem243; 
            mem244_n = (wen && ( 244 == addr))? wdata : mem244; 
            mem245_n = (wen && ( 245 == addr))? wdata : mem245; 
            mem246_n = (wen && ( 246 == addr))? wdata : mem246; 
            mem247_n = (wen && ( 247 == addr))? wdata : mem247; 
            mem248_n = (wen && ( 248 == addr))? wdata : mem248; 
            mem249_n = (wen && ( 249 == addr))? wdata : mem249; 
            mem250_n = (wen && ( 250 == addr))? wdata : mem250; 
            mem251_n = (wen && ( 251 == addr))? wdata : mem251; 
            mem252_n = (wen && ( 252 == addr))? wdata : mem252; 
            mem253_n = (wen && ( 253 == addr))? wdata : mem253; 
            mem254_n = (wen && ( 254 == addr))? wdata : mem254; 
            mem255_n = (wen && ( 255 == addr))? wdata : mem255; 
end


endmodule










